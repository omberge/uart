-- test for now...
